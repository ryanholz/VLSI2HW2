/* Parameter verilog header file */
/*
* Contains all of the parameters used throughout the design
*/

localparam L1_ADDR_WIDTH = 2;
localparam L2_ADDR_WIDTH = 3;
localparam MESI_WIDTH = 2;
localparam DATA_WIDTH = 8;
localparam NUM_CORES = 4;
localparam NUM_L1_BLOCKS = 4;
localparam NUM_L2_BLOCKS = 8;
